-- This package is used for EECS 361 from Northwestern University.
-- by Kaicheng Zhang (kaichengz@gmail.com)

library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;

package eecs361 is

  --decode
  component decode
	port(
		ins: in std_logic_vector(31 downto 0);
		regS: out std_logic_vector(4 downto 0);
		regT: out std_logic_vector(4 downto 0);
		regD: out std_logic_vector(4 downto 0);
		imm: out std_logic_vector(31 downto 0);
		opcode: out std_logic_vector(5 downto 0);
		func: out std_logic_vector(5 downto 0);
		shamt: out std_logic_vector(31 downto 0)	
	);
  end component decode;

  -- instruction
  component Instruction
	port(
		zero: in std_logic;
		clk : in std_logic;
		jump: in std_logic;
		branch: in std_logic;
		reset : in std_logic;
		instruction: out std_logic_vector(31 downto 0)		
	);
  end component Instruction;
  -- Complete_adder
  component complete_adder 
    port(
      a,b: in std_logic_vector(31 downto 0);
      ci: in std_logic;
      co,ov,zero: out std_logic;
      s: out std_logic_vector(31 downto 0)
    );
  end component complete_adder;

  -- Quarbit_adder
  component quarbit_adder
    port(
      a,b: in std_logic_vector(3 downto 0);
      ci:in std_logic;
      s:out std_logic_vector(3 downto 0);
      co,ov,zero:out std_logic
    );
  end component quarbit_adder;
  
  -- Full_Adder
  component full_adder
    port  (
      a: in std_logic;
      b: in std_logic;
      ci: in std_logic;
      s:out std_logic;
      co:out std_logic
    );
  end component full_adder;

  -- Decoders
  component dec_n
    generic (
      -- Widths of the inputs.
      n	  : integer
    );
    port (
      src   : in std_logic_vector(n-1 downto 0);
      z	    : out std_logic_vector((2**n)-1 downto 0)
    );
  end component dec_n;

  -- Multiplexors
  component mux
    port (
      sel   : in  std_logic;
      src0  : in  std_logic;
      src1  : in  std_logic;
      z     : out std_logic
    );
  end component mux;

  component mux_n
    generic (
      -- Widths of the inputs.
      n	  : integer
    );
    port (
      sel   : in  std_logic;
      src0  : in  std_logic_vector(n-1 downto 0);
      src1  : in  std_logic_vector(n-1 downto 0);
      z     : out std_logic_vector(n-1 downto 0)
    );
  end component mux_n;

  component mux_32
    port (
      sel   : in  std_logic;
      src0  : in  std_logic_vector(31 downto 0);
      src1  : in  std_logic_vector(31 downto 0);
      z	    : out std_logic_vector(31 downto 0)
    );
  end component mux_32;

  -- Flip-flops

  -- D Flip-flops from Figure C.8.4 with a falling edge trigger.
  component dff
    port (
      clk   : in  std_logic;
      d	    : in  std_logic;
      q	    : out std_logic
    );
  end component dff;

  -- D Flip-flops from Figure C.8.4 with a rising edge trigger.
  component dffr
    port (
      clk   : in  std_logic;
      d	    : in  std_logic;
      q	    : out std_logic
    );
  end component dffr;

  -- D Flip-flops from Example 13-40 in http://www.altera.com/literature/hb/qts/qts_qii51007.pdf
  component dffr_a
    port (
      clk	 : in  std_logic;
      arst   : in  std_logic;
      aload  : in  std_logic;
      adata  : in  std_logic;
      d	     : in  std_logic;
      enable : in  std_logic;
      q	     : out std_logic
    );

  end component dffr_a;

  -- A 32bit SRAM from Figure C.9.1. It can only be used for simulation.
  component sram
	generic (
	  mem_file	: string
	);
	port (
	  -- chip select
	  cs	: in  std_logic;
	  -- output enable
	  oe	: in  std_logic;
	  -- write enable
	  we	: in  std_logic;
	  -- address line
	  addr	: in  std_logic_vector(31 downto 0);
	  -- data input
	  din	: in  std_logic_vector(31 downto 0);
	  -- data output
	  dout	: out std_logic_vector(31 downto 0)
	);
  end component sram;

  -- Synchronous SRAM with asynchronous reset.
  component syncram
    generic (
	  mem_file	: string
	);
	port (
      -- clock
      clk   : in  std_logic;
	  -- chip select
	  cs	: in  std_logic;
      -- output enable
	  oe	: in  std_logic;
	  -- write enable
	  we	: in  std_logic;
	  -- address line
	  addr	: in  std_logic_vector(31 downto 0);
	  -- data input
	  din	: in  std_logic_vector(31 downto 0);
	  -- data output
	  dout	: out std_logic_vector(31 downto 0)
	);
  end component syncram;
end;
