library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;
use work.eecs361.all;

entity left_shifter is 
	port(
		a: in std_logic_vector(31 downto 0);
		s: in std_logic_vector(4 downto 0);
		result: out std_logic_vector(31 downto 0)
);
end entity left_shifter;

architecture beh of left_shifter is
signal temp0,temp1,temp2,temp3,temp4:std_logic_vector(31 downto 0);
begin
shift0_0: mux port map(src1 => '0', src0 => a(0), sel => s(0), z => temp0(0));
shift0_1: mux port map(src1 => a(0), src0 => a(1), sel => s(0), z => temp0(1));
shift0_2: mux port map(src1 => a(1), src0 => a(2), sel => s(0), z => temp0(2));
shift0_3: mux port map(src1 => a(2), src0 => a(3), sel => s(0), z => temp0(3));
shift0_4: mux port map(src1 => a(3), src0 => a(4), sel => s(0), z => temp0(4));
shift0_5: mux port map(src1 => a(4), src0 => a(5), sel => s(0), z => temp0(5));
shift0_6: mux port map(src1 => a(5), src0 => a(6), sel => s(0), z => temp0(6));
shift0_7: mux port map(src1 => a(6), src0 => a(7), sel => s(0), z => temp0(7));
shift0_8: mux port map(src1 => a(7), src0 => a(8), sel => s(0), z => temp0(8));
shift0_9: mux port map(src1 => a(8), src0 => a(9), sel => s(0), z => temp0(9));
shift0_10: mux port map(src1 => a(9), src0 => a(10), sel => s(0), z => temp0(10));
shift0_11: mux port map(src1 => a(10), src0 => a(11), sel => s(0), z => temp0(11));
shift0_12: mux port map(src1 => a(11), src0 => a(12), sel => s(0), z => temp0(12));
shift0_13: mux port map(src1 => a(12), src0 => a(13), sel => s(0), z => temp0(13));
shift0_14: mux port map(src1 => a(13), src0 => a(14), sel => s(0), z => temp0(14));
shift0_15: mux port map(src1 => a(14), src0 => a(15), sel => s(0), z => temp0(15));
shift0_16: mux port map(src1 => a(15), src0 => a(16), sel => s(0), z => temp0(16));
shift0_17: mux port map(src1 => a(16), src0 => a(17), sel => s(0), z => temp0(17));
shift0_18: mux port map(src1 => a(17), src0 => a(18), sel => s(0), z => temp0(18));
shift0_19: mux port map(src1 => a(18), src0 => a(19), sel => s(0), z => temp0(19));
shift0_20: mux port map(src1 => a(19), src0 => a(20), sel => s(0), z => temp0(20));
shift0_21: mux port map(src1 => a(20), src0 => a(21), sel => s(0), z => temp0(21));
shift0_22: mux port map(src1 => a(21), src0 => a(22), sel => s(0), z => temp0(22));
shift0_23: mux port map(src1 => a(22), src0 => a(23), sel => s(0), z => temp0(23));
shift0_24: mux port map(src1 => a(23), src0 => a(24), sel => s(0), z => temp0(24));
shift0_25: mux port map(src1 => a(24), src0 => a(25), sel => s(0), z => temp0(25));
shift0_26: mux port map(src1 => a(25), src0 => a(26), sel => s(0), z => temp0(26));
shift0_27: mux port map(src1 => a(26), src0 => a(27), sel => s(0), z => temp0(27));
shift0_28: mux port map(src1 => a(27), src0 => a(28), sel => s(0), z => temp0(28));
shift0_29: mux port map(src1 => a(28), src0 => a(29), sel => s(0), z => temp0(29));
shift0_30: mux port map(src1 => a(29), src0 => a(30), sel => s(0), z => temp0(30));
shift0_31: mux port map(src1 => a(30), src0 => a(31), sel => s(0), z => temp0(31));
shift1_0: mux port map(src1 => '0', src0 => temp0(0), sel => s(1), z => temp1(0));
shift1_1: mux port map(src1 => '0', src0 => temp0(1), sel => s(1), z => temp1(1));
shift1_2: mux port map(src1 => temp0(0), src0 => temp0(2), sel => s(1), z => temp1(2));
shift1_3: mux port map(src1 => temp0(1), src0 => temp0(3), sel => s(1), z => temp1(3));
shift1_4: mux port map(src1 => temp0(2), src0 => temp0(4), sel => s(1), z => temp1(4));
shift1_5: mux port map(src1 => temp0(3), src0 => temp0(5), sel => s(1), z => temp1(5));
shift1_6: mux port map(src1 => temp0(4), src0 => temp0(6), sel => s(1), z => temp1(6));
shift1_7: mux port map(src1 => temp0(5), src0 => temp0(7), sel => s(1), z => temp1(7));
shift1_8: mux port map(src1 => temp0(6), src0 => temp0(8), sel => s(1), z => temp1(8));
shift1_9: mux port map(src1 => temp0(7), src0 => temp0(9), sel => s(1), z => temp1(9));
shift1_10: mux port map(src1 => temp0(8), src0 => temp0(10), sel => s(1), z => temp1(10));
shift1_11: mux port map(src1 => temp0(9), src0 => temp0(11), sel => s(1), z => temp1(11));
shift1_12: mux port map(src1 => temp0(10), src0 => temp0(12), sel => s(1), z => temp1(12));
shift1_13: mux port map(src1 => temp0(11), src0 => temp0(13), sel => s(1), z => temp1(13));
shift1_14: mux port map(src1 => temp0(12), src0 => temp0(14), sel => s(1), z => temp1(14));
shift1_15: mux port map(src1 => temp0(13), src0 => temp0(15), sel => s(1), z => temp1(15));
shift1_16: mux port map(src1 => temp0(14), src0 => temp0(16), sel => s(1), z => temp1(16));
shift1_17: mux port map(src1 => temp0(15), src0 => temp0(17), sel => s(1), z => temp1(17));
shift1_18: mux port map(src1 => temp0(16), src0 => temp0(18), sel => s(1), z => temp1(18));
shift1_19: mux port map(src1 => temp0(17), src0 => temp0(19), sel => s(1), z => temp1(19));
shift1_20: mux port map(src1 => temp0(18), src0 => temp0(20), sel => s(1), z => temp1(20));
shift1_21: mux port map(src1 => temp0(19), src0 => temp0(21), sel => s(1), z => temp1(21));
shift1_22: mux port map(src1 => temp0(20), src0 => temp0(22), sel => s(1), z => temp1(22));
shift1_23: mux port map(src1 => temp0(21), src0 => temp0(23), sel => s(1), z => temp1(23));
shift1_24: mux port map(src1 => temp0(22), src0 => temp0(24), sel => s(1), z => temp1(24));
shift1_25: mux port map(src1 => temp0(23), src0 => temp0(25), sel => s(1), z => temp1(25));
shift1_26: mux port map(src1 => temp0(24), src0 => temp0(26), sel => s(1), z => temp1(26));
shift1_27: mux port map(src1 => temp0(25), src0 => temp0(27), sel => s(1), z => temp1(27));
shift1_28: mux port map(src1 => temp0(26), src0 => temp0(28), sel => s(1), z => temp1(28));
shift1_29: mux port map(src1 => temp0(27), src0 => temp0(29), sel => s(1), z => temp1(29));
shift1_30: mux port map(src1 => temp0(28), src0 => temp0(30), sel => s(1), z => temp1(30));
shift1_31: mux port map(src1 => temp0(29), src0 => temp0(31), sel => s(1), z => temp1(31));
shift2_0: mux port map(src1 => '0', src0 => temp1(0), sel => s(2), z => temp2(0));
shift2_1: mux port map(src1 => '0', src0 => temp1(1), sel => s(2), z => temp2(1));
shift2_2: mux port map(src1 => '0', src0 => temp1(2), sel => s(2), z => temp2(2));
shift2_3: mux port map(src1 => '0', src0 => temp1(3), sel => s(2), z => temp2(3));
shift2_4: mux port map(src1 => temp1(0), src0 => temp1(4), sel => s(2), z => temp2(4));
shift2_5: mux port map(src1 => temp1(1), src0 => temp1(5), sel => s(2), z => temp2(5));
shift2_6: mux port map(src1 => temp1(2), src0 => temp1(6), sel => s(2), z => temp2(6));
shift2_7: mux port map(src1 => temp1(3), src0 => temp1(7), sel => s(2), z => temp2(7));
shift2_8: mux port map(src1 => temp1(4), src0 => temp1(8), sel => s(2), z => temp2(8));
shift2_9: mux port map(src1 => temp1(5), src0 => temp1(9), sel => s(2), z => temp2(9));
shift2_10: mux port map(src1 => temp1(6), src0 => temp1(10), sel => s(2), z => temp2(10));
shift2_11: mux port map(src1 => temp1(7), src0 => temp1(11), sel => s(2), z => temp2(11));
shift2_12: mux port map(src1 => temp1(8), src0 => temp1(12), sel => s(2), z => temp2(12));
shift2_13: mux port map(src1 => temp1(9), src0 => temp1(13), sel => s(2), z => temp2(13));
shift2_14: mux port map(src1 => temp1(10), src0 => temp1(14), sel => s(2), z => temp2(14));
shift2_15: mux port map(src1 => temp1(11), src0 => temp1(15), sel => s(2), z => temp2(15));
shift2_16: mux port map(src1 => temp1(12), src0 => temp1(16), sel => s(2), z => temp2(16));
shift2_17: mux port map(src1 => temp1(13), src0 => temp1(17), sel => s(2), z => temp2(17));
shift2_18: mux port map(src1 => temp1(14), src0 => temp1(18), sel => s(2), z => temp2(18));
shift2_19: mux port map(src1 => temp1(15), src0 => temp1(19), sel => s(2), z => temp2(19));
shift2_20: mux port map(src1 => temp1(16), src0 => temp1(20), sel => s(2), z => temp2(20));
shift2_21: mux port map(src1 => temp1(17), src0 => temp1(21), sel => s(2), z => temp2(21));
shift2_22: mux port map(src1 => temp1(18), src0 => temp1(22), sel => s(2), z => temp2(22));
shift2_23: mux port map(src1 => temp1(19), src0 => temp1(23), sel => s(2), z => temp2(23));
shift2_24: mux port map(src1 => temp1(20), src0 => temp1(24), sel => s(2), z => temp2(24));
shift2_25: mux port map(src1 => temp1(21), src0 => temp1(25), sel => s(2), z => temp2(25));
shift2_26: mux port map(src1 => temp1(22), src0 => temp1(26), sel => s(2), z => temp2(26));
shift2_27: mux port map(src1 => temp1(23), src0 => temp1(27), sel => s(2), z => temp2(27));
shift2_28: mux port map(src1 => temp1(24), src0 => temp1(28), sel => s(2), z => temp2(28));
shift2_29: mux port map(src1 => temp1(25), src0 => temp1(29), sel => s(2), z => temp2(29));
shift2_30: mux port map(src1 => temp1(26), src0 => temp1(30), sel => s(2), z => temp2(30));
shift2_31: mux port map(src1 => temp1(27), src0 => temp1(31), sel => s(2), z => temp2(31));
shift3_0: mux port map(src1 => '0', src0 => temp2(0), sel => s(3), z => temp3(0));
shift3_1: mux port map(src1 => '0', src0 => temp2(1), sel => s(3), z => temp3(1));
shift3_2: mux port map(src1 => '0', src0 => temp2(2), sel => s(3), z => temp3(2));
shift3_3: mux port map(src1 => '0', src0 => temp2(3), sel => s(3), z => temp3(3));
shift3_4: mux port map(src1 => '0', src0 => temp2(4), sel => s(3), z => temp3(4));
shift3_5: mux port map(src1 => '0', src0 => temp2(5), sel => s(3), z => temp3(5));
shift3_6: mux port map(src1 => '0', src0 => temp2(6), sel => s(3), z => temp3(6));
shift3_7: mux port map(src1 => '0', src0 => temp2(7), sel => s(3), z => temp3(7));
shift3_8: mux port map(src1 => temp2(0), src0 => temp2(8), sel => s(3), z => temp3(8));
shift3_9: mux port map(src1 => temp2(1), src0 => temp2(9), sel => s(3), z => temp3(9));
shift3_10: mux port map(src1 => temp2(2), src0 => temp2(10), sel => s(3), z => temp3(10));
shift3_11: mux port map(src1 => temp2(3), src0 => temp2(11), sel => s(3), z => temp3(11));
shift3_12: mux port map(src1 => temp2(4), src0 => temp2(12), sel => s(3), z => temp3(12));
shift3_13: mux port map(src1 => temp2(5), src0 => temp2(13), sel => s(3), z => temp3(13));
shift3_14: mux port map(src1 => temp2(6), src0 => temp2(14), sel => s(3), z => temp3(14));
shift3_15: mux port map(src1 => temp2(7), src0 => temp2(15), sel => s(3), z => temp3(15));
shift3_16: mux port map(src1 => temp2(8), src0 => temp2(16), sel => s(3), z => temp3(16));
shift3_17: mux port map(src1 => temp2(9), src0 => temp2(17), sel => s(3), z => temp3(17));
shift3_18: mux port map(src1 => temp2(10), src0 => temp2(18), sel => s(3), z => temp3(18));
shift3_19: mux port map(src1 => temp2(11), src0 => temp2(19), sel => s(3), z => temp3(19));
shift3_20: mux port map(src1 => temp2(12), src0 => temp2(20), sel => s(3), z => temp3(20));
shift3_21: mux port map(src1 => temp2(13), src0 => temp2(21), sel => s(3), z => temp3(21));
shift3_22: mux port map(src1 => temp2(14), src0 => temp2(22), sel => s(3), z => temp3(22));
shift3_23: mux port map(src1 => temp2(15), src0 => temp2(23), sel => s(3), z => temp3(23));
shift3_24: mux port map(src1 => temp2(16), src0 => temp2(24), sel => s(3), z => temp3(24));
shift3_25: mux port map(src1 => temp2(17), src0 => temp2(25), sel => s(3), z => temp3(25));
shift3_26: mux port map(src1 => temp2(18), src0 => temp2(26), sel => s(3), z => temp3(26));
shift3_27: mux port map(src1 => temp2(19), src0 => temp2(27), sel => s(3), z => temp3(27));
shift3_28: mux port map(src1 => temp2(20), src0 => temp2(28), sel => s(3), z => temp3(28));
shift3_29: mux port map(src1 => temp2(21), src0 => temp2(29), sel => s(3), z => temp3(29));
shift3_30: mux port map(src1 => temp2(22), src0 => temp2(30), sel => s(3), z => temp3(30));
shift3_31: mux port map(src1 => temp2(23), src0 => temp2(31), sel => s(3), z => temp3(31));
shift4_0: mux port map(src1 => '0', src0 => temp3(0), sel => s(4), z => temp4(0));
shift4_1: mux port map(src1 => '0', src0 => temp3(1), sel => s(4), z => temp4(1));
shift4_2: mux port map(src1 => '0', src0 => temp3(2), sel => s(4), z => temp4(2));
shift4_3: mux port map(src1 => '0', src0 => temp3(3), sel => s(4), z => temp4(3));
shift4_4: mux port map(src1 => '0', src0 => temp3(4), sel => s(4), z => temp4(4));
shift4_5: mux port map(src1 => '0', src0 => temp3(5), sel => s(4), z => temp4(5));
shift4_6: mux port map(src1 => '0', src0 => temp3(6), sel => s(4), z => temp4(6));
shift4_7: mux port map(src1 => '0', src0 => temp3(7), sel => s(4), z => temp4(7));
shift4_8: mux port map(src1 => '0', src0 => temp3(8), sel => s(4), z => temp4(8));
shift4_9: mux port map(src1 => '0', src0 => temp3(9), sel => s(4), z => temp4(9));
shift4_10: mux port map(src1 => '0', src0 => temp3(10), sel => s(4), z => temp4(10));
shift4_11: mux port map(src1 => '0', src0 => temp3(11), sel => s(4), z => temp4(11));
shift4_12: mux port map(src1 => '0', src0 => temp3(12), sel => s(4), z => temp4(12));
shift4_13: mux port map(src1 => '0', src0 => temp3(13), sel => s(4), z => temp4(13));
shift4_14: mux port map(src1 => '0', src0 => temp3(14), sel => s(4), z => temp4(14));
shift4_15: mux port map(src1 => '0', src0 => temp3(15), sel => s(4), z => temp4(15));
shift4_16: mux port map(src1 => temp3(0), src0 => temp3(16), sel => s(4), z => temp4(16));
shift4_17: mux port map(src1 => temp3(1), src0 => temp3(17), sel => s(4), z => temp4(17));
shift4_18: mux port map(src1 => temp3(2), src0 => temp3(18), sel => s(4), z => temp4(18));
shift4_19: mux port map(src1 => temp3(3), src0 => temp3(19), sel => s(4), z => temp4(19));
shift4_20: mux port map(src1 => temp3(4), src0 => temp3(20), sel => s(4), z => temp4(20));
shift4_21: mux port map(src1 => temp3(5), src0 => temp3(21), sel => s(4), z => temp4(21));
shift4_22: mux port map(src1 => temp3(6), src0 => temp3(22), sel => s(4), z => temp4(22));
shift4_23: mux port map(src1 => temp3(7), src0 => temp3(23), sel => s(4), z => temp4(23));
shift4_24: mux port map(src1 => temp3(8), src0 => temp3(24), sel => s(4), z => temp4(24));
shift4_25: mux port map(src1 => temp3(9), src0 => temp3(25), sel => s(4), z => temp4(25));
shift4_26: mux port map(src1 => temp3(10), src0 => temp3(26), sel => s(4), z => temp4(26));
shift4_27: mux port map(src1 => temp3(11), src0 => temp3(27), sel => s(4), z => temp4(27));
shift4_28: mux port map(src1 => temp3(12), src0 => temp3(28), sel => s(4), z => temp4(28));
shift4_29: mux port map(src1 => temp3(13), src0 => temp3(29), sel => s(4), z => temp4(29));
shift4_30: mux port map(src1 => temp3(14), src0 => temp3(30), sel => s(4), z => temp4(30));
shift4_31: mux port map(src1 => temp3(15), src0 => temp3(31), sel => s(4), z => temp4(31));
result <= temp4;
end beh;
